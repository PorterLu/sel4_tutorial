arch x86_64

objects {
cnode_client_1 = cnode (3 bits)
cnode_client_2 = cnode (3 bits)
cnode_server = cnode (3 bits)
endpoint = ep
frame_client_1_0000 = frame (4k, fill: [{0 548 CDL_FrameFill_FileData "client_1" 0}])
frame_client_1_0001 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_1" 4096}])
frame_client_1_0002 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_1" 8192}])
frame_client_1_0003 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_1" 12288}])
frame_client_1_0004 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_1" 16384}])
frame_client_1_0005 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_1" 20480}])
frame_client_1_0006 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_1" 24576}])
frame_client_1_0007 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_1" 28672}])
frame_client_1_0008 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_1" 32768}])
frame_client_1_0009 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_1" 36864}])
frame_client_1_0010 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_1" 40960}])
frame_client_1_0011 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_1" 45056}])
frame_client_1_0012 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_1" 49152}])
frame_client_1_0013 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_1" 53248}])
frame_client_1_0014 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_1" 57344}])
frame_client_1_0015 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_1" 61440}])
frame_client_1_0016 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_1" 65536}])
frame_client_1_0017 = frame (4k, fill: [{0 2207 CDL_FrameFill_FileData "client_1" 69632}])
frame_client_1_0018 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_1" 73728}])
frame_client_1_0019 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_1" 77824}])
frame_client_1_0020 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_1" 81920}])
frame_client_1_0021 = frame (4k, fill: [{0 2800 CDL_FrameFill_FileData "client_1" 86016}])
frame_client_1_0022 = frame (4k, fill: [{4040 56 CDL_FrameFill_FileData "client_1" 90056}])
frame_client_1_0023 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_1" 90112}])
frame_client_1_0024 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_1" 94208}])
frame_client_1_0042 = frame (4k, fill: [{0 8 CDL_FrameFill_FileData "client_1" 167936}])
frame_client_1_0043 = frame (4k, fill: [])
frame_client_1_0044 = frame (4k, fill: [])
frame_client_1_0045 = frame (4k, fill: [])
frame_client_1_0046 = frame (4k, fill: [])
frame_client_1_0047 = frame (4k, fill: [])
frame_client_1_0048 = frame (4k, fill: [])
frame_client_1_0049 = frame (4k, fill: [])
frame_client_1_0050 = frame (4k, fill: [])
frame_client_1_0051 = frame (4k, fill: [])
frame_client_1_0052 = frame (4k, fill: [])
frame_client_1_0053 = frame (4k, fill: [])
frame_client_1_0054 = frame (4k, fill: [])
frame_client_1_0055 = frame (4k, fill: [])
frame_client_1_0056 = frame (4k, fill: [])
frame_client_1_0057 = frame (4k, fill: [])
frame_client_1_0058 = frame (4k, fill: [])
frame_client_1_0059 = frame (4k, fill: [])
frame_client_1_0060 = frame (4k, fill: [])
frame_client_1_0061 = frame (4k, fill: [])
frame_client_1_0062 = frame (4k, fill: [])
frame_client_1_0063 = frame (4k, fill: [])
frame_client_1_0064 = frame (4k, fill: [])
frame_client_1_0065 = frame (4k, fill: [])
frame_client_1_0066 = frame (4k, fill: [])
frame_client_1_0067 = frame (4k, fill: [])
frame_client_1_0068 = frame (4k, fill: [])
frame_client_1_0069 = frame (4k, fill: [])
frame_client_1_0070 = frame (4k, fill: [])
frame_client_1_0071 = frame (4k, fill: [])
frame_client_1_0072 = frame (4k, fill: [])
frame_client_1_0073 = frame (4k, fill: [])
frame_client_1_0074 = frame (4k, fill: [])
frame_client_1_0075 = frame (4k, fill: [])
frame_client_1_0076 = frame (4k, fill: [])
frame_client_1_0077 = frame (4k, fill: [])
frame_client_1_0078 = frame (4k, fill: [])
frame_client_1_0079 = frame (4k, fill: [])
frame_client_1_0080 = frame (4k, fill: [])
frame_client_1_0081 = frame (4k, fill: [])
frame_client_1_0082 = frame (4k, fill: [])
frame_client_1_0083 = frame (4k, fill: [])
frame_client_1_0084 = frame (4k, fill: [])
frame_client_1_0085 = frame (4k, fill: [])
frame_client_1_0086 = frame (4k, fill: [])
frame_client_1_0087 = frame (4k, fill: [])
frame_client_1_0088 = frame (4k, fill: [])
frame_client_1_0089 = frame (4k, fill: [])
frame_client_1_0090 = frame (4k, fill: [])
frame_client_1_0091 = frame (4k, fill: [])
frame_client_1_0092 = frame (4k, fill: [])
frame_client_1_0093 = frame (4k, fill: [])
frame_client_1_0094 = frame (4k, fill: [])
frame_client_1_0095 = frame (4k, fill: [])
frame_client_1_0096 = frame (4k, fill: [])
frame_client_1_0097 = frame (4k, fill: [])
frame_client_1_0098 = frame (4k, fill: [])
frame_client_1_0099 = frame (4k, fill: [])
frame_client_1_0100 = frame (4k, fill: [])
frame_client_1_0101 = frame (4k, fill: [])
frame_client_1_0102 = frame (4k, fill: [])
frame_client_1_0103 = frame (4k, fill: [])
frame_client_1_0104 = frame (4k, fill: [])
frame_client_1_0105 = frame (4k, fill: [])
frame_client_1_0106 = frame (4k, fill: [])
frame_client_1_0107 = frame (4k, fill: [])
frame_client_1_0108 = frame (4k, fill: [])
frame_client_1_0109 = frame (4k, fill: [])
frame_client_1_0110 = frame (4k, fill: [])
frame_client_1_0111 = frame (4k, fill: [])
frame_client_1_0112 = frame (4k, fill: [])
frame_client_1_0113 = frame (4k, fill: [])
frame_client_1_0114 = frame (4k, fill: [])
frame_client_1_0115 = frame (4k, fill: [])
frame_client_1_0116 = frame (4k, fill: [])
frame_client_1_0117 = frame (4k, fill: [])
frame_client_1_0118 = frame (4k, fill: [])
frame_client_1_0119 = frame (4k, fill: [])
frame_client_1_0120 = frame (4k, fill: [])
frame_client_1_0121 = frame (4k, fill: [])
frame_client_1_0122 = frame (4k, fill: [])
frame_client_1_0123 = frame (4k, fill: [])
frame_client_1_0124 = frame (4k, fill: [])
frame_client_1_0125 = frame (4k, fill: [])
frame_client_1_0126 = frame (4k, fill: [])
frame_client_1_0127 = frame (4k, fill: [])
frame_client_1_0128 = frame (4k, fill: [])
frame_client_1_0129 = frame (4k, fill: [])
frame_client_1_0130 = frame (4k, fill: [])
frame_client_1_0131 = frame (4k, fill: [])
frame_client_1_0132 = frame (4k, fill: [])
frame_client_1_0133 = frame (4k, fill: [])
frame_client_1_0134 = frame (4k, fill: [])
frame_client_1_0135 = frame (4k, fill: [])
frame_client_1_0136 = frame (4k, fill: [])
frame_client_1_0137 = frame (4k, fill: [])
frame_client_1_0138 = frame (4k, fill: [])
frame_client_1_0139 = frame (4k, fill: [])
frame_client_1_0140 = frame (4k, fill: [])
frame_client_1_0141 = frame (4k, fill: [])
frame_client_1_0142 = frame (4k, fill: [])
frame_client_1_0143 = frame (4k, fill: [])
frame_client_1_0144 = frame (4k, fill: [])
frame_client_1_0145 = frame (4k, fill: [])
frame_client_1_0146 = frame (4k, fill: [])
frame_client_1_0147 = frame (4k, fill: [])
frame_client_1_0148 = frame (4k, fill: [])
frame_client_1_0149 = frame (4k, fill: [])
frame_client_1_0150 = frame (4k, fill: [])
frame_client_1_0151 = frame (4k, fill: [])
frame_client_1_0152 = frame (4k, fill: [])
frame_client_1_0153 = frame (4k, fill: [])
frame_client_1_0154 = frame (4k, fill: [])
frame_client_1_0155 = frame (4k, fill: [])
frame_client_1_0156 = frame (4k, fill: [])
frame_client_1_0157 = frame (4k, fill: [])
frame_client_1_0158 = frame (4k, fill: [])
frame_client_1_0159 = frame (4k, fill: [])
frame_client_1_0160 = frame (4k, fill: [])
frame_client_1_0161 = frame (4k, fill: [])
frame_client_1_0162 = frame (4k, fill: [])
frame_client_1_0163 = frame (4k, fill: [])
frame_client_1_0164 = frame (4k, fill: [])
frame_client_1_0165 = frame (4k, fill: [])
frame_client_1_0166 = frame (4k, fill: [])
frame_client_1_0167 = frame (4k, fill: [])
frame_client_1_0168 = frame (4k, fill: [])
frame_client_1_0169 = frame (4k, fill: [])
frame_client_1_0170 = frame (4k, fill: [])
frame_client_1_0171 = frame (4k, fill: [])
frame_client_1_0172 = frame (4k, fill: [])
frame_client_1_0173 = frame (4k, fill: [])
frame_client_1_0174 = frame (4k, fill: [])
frame_client_1_0175 = frame (4k, fill: [])
frame_client_1_0176 = frame (4k, fill: [])
frame_client_1_0177 = frame (4k, fill: [])
frame_client_1_0178 = frame (4k, fill: [])
frame_client_1_0179 = frame (4k, fill: [])
frame_client_1_0180 = frame (4k, fill: [])
frame_client_1_0181 = frame (4k, fill: [])
frame_client_1_0182 = frame (4k, fill: [])
frame_client_1_0183 = frame (4k, fill: [])
frame_client_1_0184 = frame (4k, fill: [])
frame_client_1_0185 = frame (4k, fill: [])
frame_client_1_0186 = frame (4k, fill: [])
frame_client_1_0187 = frame (4k, fill: [])
frame_client_1_0188 = frame (4k, fill: [])
frame_client_1_0189 = frame (4k, fill: [])
frame_client_1_0190 = frame (4k, fill: [])
frame_client_1_0191 = frame (4k, fill: [])
frame_client_1_0192 = frame (4k, fill: [])
frame_client_1_0193 = frame (4k, fill: [])
frame_client_1_0194 = frame (4k, fill: [])
frame_client_1_0195 = frame (4k, fill: [])
frame_client_1_0196 = frame (4k, fill: [])
frame_client_1_0197 = frame (4k, fill: [])
frame_client_1_0198 = frame (4k, fill: [])
frame_client_1_0199 = frame (4k, fill: [])
frame_client_1_0200 = frame (4k, fill: [])
frame_client_1_0201 = frame (4k, fill: [])
frame_client_1_0202 = frame (4k, fill: [])
frame_client_1_0203 = frame (4k, fill: [])
frame_client_1_0204 = frame (4k, fill: [])
frame_client_1_0205 = frame (4k, fill: [])
frame_client_1_0206 = frame (4k, fill: [])
frame_client_1_0207 = frame (4k, fill: [])
frame_client_1_0208 = frame (4k, fill: [])
frame_client_1_0209 = frame (4k, fill: [])
frame_client_1_0210 = frame (4k, fill: [])
frame_client_1_0211 = frame (4k, fill: [])
frame_client_1_0212 = frame (4k, fill: [])
frame_client_1_0213 = frame (4k, fill: [])
frame_client_1_0214 = frame (4k, fill: [])
frame_client_1_0215 = frame (4k, fill: [])
frame_client_1_0216 = frame (4k, fill: [])
frame_client_1_0217 = frame (4k, fill: [])
frame_client_1_0218 = frame (4k, fill: [])
frame_client_1_0219 = frame (4k, fill: [])
frame_client_1_0220 = frame (4k, fill: [])
frame_client_1_0221 = frame (4k, fill: [])
frame_client_1_0222 = frame (4k, fill: [])
frame_client_1_0223 = frame (4k, fill: [])
frame_client_1_0224 = frame (4k, fill: [])
frame_client_1_0225 = frame (4k, fill: [])
frame_client_1_0226 = frame (4k, fill: [])
frame_client_1_0227 = frame (4k, fill: [])
frame_client_1_0228 = frame (4k, fill: [])
frame_client_1_0229 = frame (4k, fill: [])
frame_client_1_0230 = frame (4k, fill: [])
frame_client_1_0231 = frame (4k, fill: [])
frame_client_1_0232 = frame (4k, fill: [])
frame_client_1_0233 = frame (4k, fill: [])
frame_client_1_0234 = frame (4k, fill: [])
frame_client_1_0235 = frame (4k, fill: [])
frame_client_1_0236 = frame (4k, fill: [])
frame_client_1_0237 = frame (4k, fill: [])
frame_client_1_0238 = frame (4k, fill: [])
frame_client_1_0239 = frame (4k, fill: [])
frame_client_1_0240 = frame (4k, fill: [])
frame_client_1_0241 = frame (4k, fill: [])
frame_client_1_0242 = frame (4k, fill: [])
frame_client_1_0243 = frame (4k, fill: [])
frame_client_1_0244 = frame (4k, fill: [])
frame_client_1_0245 = frame (4k, fill: [])
frame_client_1_0246 = frame (4k, fill: [])
frame_client_1_0247 = frame (4k, fill: [])
frame_client_1_0248 = frame (4k, fill: [])
frame_client_1_0249 = frame (4k, fill: [])
frame_client_1_0250 = frame (4k, fill: [])
frame_client_1_0251 = frame (4k, fill: [])
frame_client_1_0252 = frame (4k, fill: [])
frame_client_1_0253 = frame (4k, fill: [])
frame_client_1_0254 = frame (4k, fill: [])
frame_client_1_0255 = frame (4k, fill: [])
frame_client_1_0256 = frame (4k, fill: [])
frame_client_1_0257 = frame (4k, fill: [])
frame_client_1_0258 = frame (4k, fill: [])
frame_client_1_0259 = frame (4k, fill: [])
frame_client_1_0260 = frame (4k, fill: [])
frame_client_1_0261 = frame (4k, fill: [])
frame_client_1_0262 = frame (4k, fill: [])
frame_client_1_0263 = frame (4k, fill: [])
frame_client_1_0264 = frame (4k, fill: [])
frame_client_1_0265 = frame (4k, fill: [])
frame_client_1_0266 = frame (4k, fill: [])
frame_client_1_0267 = frame (4k, fill: [])
frame_client_1_0268 = frame (4k, fill: [])
frame_client_1_0269 = frame (4k, fill: [])
frame_client_1_0270 = frame (4k, fill: [])
frame_client_1_0271 = frame (4k, fill: [])
frame_client_1_0272 = frame (4k, fill: [])
frame_client_1_0273 = frame (4k, fill: [])
frame_client_1_0274 = frame (4k, fill: [])
frame_client_1_0275 = frame (4k, fill: [])
frame_client_1_0276 = frame (4k, fill: [])
frame_client_1_0277 = frame (4k, fill: [])
frame_client_1_0278 = frame (4k, fill: [])
frame_client_1_0279 = frame (4k, fill: [])
frame_client_1_0280 = frame (4k, fill: [])
frame_client_1_0281 = frame (4k, fill: [])
frame_client_1_0282 = frame (4k, fill: [])
frame_client_1_0283 = frame (4k, fill: [])
frame_client_1_0284 = frame (4k, fill: [])
frame_client_1_0285 = frame (4k, fill: [])
frame_client_1_0286 = frame (4k, fill: [])
frame_client_1_0287 = frame (4k, fill: [])
frame_client_1_0288 = frame (4k, fill: [])
frame_client_1_0289 = frame (4k, fill: [])
frame_client_1_0290 = frame (4k, fill: [])
frame_client_1_0291 = frame (4k, fill: [])
frame_client_1_0292 = frame (4k, fill: [])
frame_client_1_0293 = frame (4k, fill: [])
frame_client_1_0294 = frame (4k, fill: [])
frame_client_1_0295 = frame (4k, fill: [])
frame_client_1_0296 = frame (4k, fill: [])
frame_client_1_0297 = frame (4k, fill: [])
frame_client_1_0298 = frame (4k, fill: [])
frame_client_1_0299 = frame (4k, fill: [])
frame_client_1_0300 = frame (4k, fill: [])
frame_client_1_0301 = frame (4k, fill: [])
frame_client_1_0302 = frame (4k, fill: [])
frame_client_1_0303 = frame (4k, fill: [])
frame_client_1_0304 = frame (4k, fill: [])
frame_client_1_0305 = frame (4k, fill: [])
frame_client_2_0000 = frame (4k, fill: [{0 548 CDL_FrameFill_FileData "client_2" 0}])
frame_client_2_0001 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_2" 4096}])
frame_client_2_0002 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_2" 8192}])
frame_client_2_0003 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_2" 12288}])
frame_client_2_0004 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_2" 16384}])
frame_client_2_0005 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_2" 20480}])
frame_client_2_0006 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_2" 24576}])
frame_client_2_0007 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_2" 28672}])
frame_client_2_0008 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_2" 32768}])
frame_client_2_0009 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_2" 36864}])
frame_client_2_0010 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_2" 40960}])
frame_client_2_0011 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_2" 45056}])
frame_client_2_0012 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_2" 49152}])
frame_client_2_0013 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_2" 53248}])
frame_client_2_0014 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_2" 57344}])
frame_client_2_0015 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_2" 61440}])
frame_client_2_0016 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_2" 65536}])
frame_client_2_0017 = frame (4k, fill: [{0 2207 CDL_FrameFill_FileData "client_2" 69632}])
frame_client_2_0018 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_2" 73728}])
frame_client_2_0019 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_2" 77824}])
frame_client_2_0020 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_2" 81920}])
frame_client_2_0021 = frame (4k, fill: [{0 2800 CDL_FrameFill_FileData "client_2" 86016}])
frame_client_2_0022 = frame (4k, fill: [{4040 56 CDL_FrameFill_FileData "client_2" 90056}])
frame_client_2_0023 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_2" 90112}])
frame_client_2_0024 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_2" 94208}])
frame_client_2_0042 = frame (4k, fill: [{0 8 CDL_FrameFill_FileData "client_2" 167936}])
frame_client_2_0043 = frame (4k, fill: [])
frame_client_2_0044 = frame (4k, fill: [])
frame_client_2_0045 = frame (4k, fill: [])
frame_client_2_0046 = frame (4k, fill: [])
frame_client_2_0047 = frame (4k, fill: [])
frame_client_2_0048 = frame (4k, fill: [])
frame_client_2_0049 = frame (4k, fill: [])
frame_client_2_0050 = frame (4k, fill: [])
frame_client_2_0051 = frame (4k, fill: [])
frame_client_2_0052 = frame (4k, fill: [])
frame_client_2_0053 = frame (4k, fill: [])
frame_client_2_0054 = frame (4k, fill: [])
frame_client_2_0055 = frame (4k, fill: [])
frame_client_2_0056 = frame (4k, fill: [])
frame_client_2_0057 = frame (4k, fill: [])
frame_client_2_0058 = frame (4k, fill: [])
frame_client_2_0059 = frame (4k, fill: [])
frame_client_2_0060 = frame (4k, fill: [])
frame_client_2_0061 = frame (4k, fill: [])
frame_client_2_0062 = frame (4k, fill: [])
frame_client_2_0063 = frame (4k, fill: [])
frame_client_2_0064 = frame (4k, fill: [])
frame_client_2_0065 = frame (4k, fill: [])
frame_client_2_0066 = frame (4k, fill: [])
frame_client_2_0067 = frame (4k, fill: [])
frame_client_2_0068 = frame (4k, fill: [])
frame_client_2_0069 = frame (4k, fill: [])
frame_client_2_0070 = frame (4k, fill: [])
frame_client_2_0071 = frame (4k, fill: [])
frame_client_2_0072 = frame (4k, fill: [])
frame_client_2_0073 = frame (4k, fill: [])
frame_client_2_0074 = frame (4k, fill: [])
frame_client_2_0075 = frame (4k, fill: [])
frame_client_2_0076 = frame (4k, fill: [])
frame_client_2_0077 = frame (4k, fill: [])
frame_client_2_0078 = frame (4k, fill: [])
frame_client_2_0079 = frame (4k, fill: [])
frame_client_2_0080 = frame (4k, fill: [])
frame_client_2_0081 = frame (4k, fill: [])
frame_client_2_0082 = frame (4k, fill: [])
frame_client_2_0083 = frame (4k, fill: [])
frame_client_2_0084 = frame (4k, fill: [])
frame_client_2_0085 = frame (4k, fill: [])
frame_client_2_0086 = frame (4k, fill: [])
frame_client_2_0087 = frame (4k, fill: [])
frame_client_2_0088 = frame (4k, fill: [])
frame_client_2_0089 = frame (4k, fill: [])
frame_client_2_0090 = frame (4k, fill: [])
frame_client_2_0091 = frame (4k, fill: [])
frame_client_2_0092 = frame (4k, fill: [])
frame_client_2_0093 = frame (4k, fill: [])
frame_client_2_0094 = frame (4k, fill: [])
frame_client_2_0095 = frame (4k, fill: [])
frame_client_2_0096 = frame (4k, fill: [])
frame_client_2_0097 = frame (4k, fill: [])
frame_client_2_0098 = frame (4k, fill: [])
frame_client_2_0099 = frame (4k, fill: [])
frame_client_2_0100 = frame (4k, fill: [])
frame_client_2_0101 = frame (4k, fill: [])
frame_client_2_0102 = frame (4k, fill: [])
frame_client_2_0103 = frame (4k, fill: [])
frame_client_2_0104 = frame (4k, fill: [])
frame_client_2_0105 = frame (4k, fill: [])
frame_client_2_0106 = frame (4k, fill: [])
frame_client_2_0107 = frame (4k, fill: [])
frame_client_2_0108 = frame (4k, fill: [])
frame_client_2_0109 = frame (4k, fill: [])
frame_client_2_0110 = frame (4k, fill: [])
frame_client_2_0111 = frame (4k, fill: [])
frame_client_2_0112 = frame (4k, fill: [])
frame_client_2_0113 = frame (4k, fill: [])
frame_client_2_0114 = frame (4k, fill: [])
frame_client_2_0115 = frame (4k, fill: [])
frame_client_2_0116 = frame (4k, fill: [])
frame_client_2_0117 = frame (4k, fill: [])
frame_client_2_0118 = frame (4k, fill: [])
frame_client_2_0119 = frame (4k, fill: [])
frame_client_2_0120 = frame (4k, fill: [])
frame_client_2_0121 = frame (4k, fill: [])
frame_client_2_0122 = frame (4k, fill: [])
frame_client_2_0123 = frame (4k, fill: [])
frame_client_2_0124 = frame (4k, fill: [])
frame_client_2_0125 = frame (4k, fill: [])
frame_client_2_0126 = frame (4k, fill: [])
frame_client_2_0127 = frame (4k, fill: [])
frame_client_2_0128 = frame (4k, fill: [])
frame_client_2_0129 = frame (4k, fill: [])
frame_client_2_0130 = frame (4k, fill: [])
frame_client_2_0131 = frame (4k, fill: [])
frame_client_2_0132 = frame (4k, fill: [])
frame_client_2_0133 = frame (4k, fill: [])
frame_client_2_0134 = frame (4k, fill: [])
frame_client_2_0135 = frame (4k, fill: [])
frame_client_2_0136 = frame (4k, fill: [])
frame_client_2_0137 = frame (4k, fill: [])
frame_client_2_0138 = frame (4k, fill: [])
frame_client_2_0139 = frame (4k, fill: [])
frame_client_2_0140 = frame (4k, fill: [])
frame_client_2_0141 = frame (4k, fill: [])
frame_client_2_0142 = frame (4k, fill: [])
frame_client_2_0143 = frame (4k, fill: [])
frame_client_2_0144 = frame (4k, fill: [])
frame_client_2_0145 = frame (4k, fill: [])
frame_client_2_0146 = frame (4k, fill: [])
frame_client_2_0147 = frame (4k, fill: [])
frame_client_2_0148 = frame (4k, fill: [])
frame_client_2_0149 = frame (4k, fill: [])
frame_client_2_0150 = frame (4k, fill: [])
frame_client_2_0151 = frame (4k, fill: [])
frame_client_2_0152 = frame (4k, fill: [])
frame_client_2_0153 = frame (4k, fill: [])
frame_client_2_0154 = frame (4k, fill: [])
frame_client_2_0155 = frame (4k, fill: [])
frame_client_2_0156 = frame (4k, fill: [])
frame_client_2_0157 = frame (4k, fill: [])
frame_client_2_0158 = frame (4k, fill: [])
frame_client_2_0159 = frame (4k, fill: [])
frame_client_2_0160 = frame (4k, fill: [])
frame_client_2_0161 = frame (4k, fill: [])
frame_client_2_0162 = frame (4k, fill: [])
frame_client_2_0163 = frame (4k, fill: [])
frame_client_2_0164 = frame (4k, fill: [])
frame_client_2_0165 = frame (4k, fill: [])
frame_client_2_0166 = frame (4k, fill: [])
frame_client_2_0167 = frame (4k, fill: [])
frame_client_2_0168 = frame (4k, fill: [])
frame_client_2_0169 = frame (4k, fill: [])
frame_client_2_0170 = frame (4k, fill: [])
frame_client_2_0171 = frame (4k, fill: [])
frame_client_2_0172 = frame (4k, fill: [])
frame_client_2_0173 = frame (4k, fill: [])
frame_client_2_0174 = frame (4k, fill: [])
frame_client_2_0175 = frame (4k, fill: [])
frame_client_2_0176 = frame (4k, fill: [])
frame_client_2_0177 = frame (4k, fill: [])
frame_client_2_0178 = frame (4k, fill: [])
frame_client_2_0179 = frame (4k, fill: [])
frame_client_2_0180 = frame (4k, fill: [])
frame_client_2_0181 = frame (4k, fill: [])
frame_client_2_0182 = frame (4k, fill: [])
frame_client_2_0183 = frame (4k, fill: [])
frame_client_2_0184 = frame (4k, fill: [])
frame_client_2_0185 = frame (4k, fill: [])
frame_client_2_0186 = frame (4k, fill: [])
frame_client_2_0187 = frame (4k, fill: [])
frame_client_2_0188 = frame (4k, fill: [])
frame_client_2_0189 = frame (4k, fill: [])
frame_client_2_0190 = frame (4k, fill: [])
frame_client_2_0191 = frame (4k, fill: [])
frame_client_2_0192 = frame (4k, fill: [])
frame_client_2_0193 = frame (4k, fill: [])
frame_client_2_0194 = frame (4k, fill: [])
frame_client_2_0195 = frame (4k, fill: [])
frame_client_2_0196 = frame (4k, fill: [])
frame_client_2_0197 = frame (4k, fill: [])
frame_client_2_0198 = frame (4k, fill: [])
frame_client_2_0199 = frame (4k, fill: [])
frame_client_2_0200 = frame (4k, fill: [])
frame_client_2_0201 = frame (4k, fill: [])
frame_client_2_0202 = frame (4k, fill: [])
frame_client_2_0203 = frame (4k, fill: [])
frame_client_2_0204 = frame (4k, fill: [])
frame_client_2_0205 = frame (4k, fill: [])
frame_client_2_0206 = frame (4k, fill: [])
frame_client_2_0207 = frame (4k, fill: [])
frame_client_2_0208 = frame (4k, fill: [])
frame_client_2_0209 = frame (4k, fill: [])
frame_client_2_0210 = frame (4k, fill: [])
frame_client_2_0211 = frame (4k, fill: [])
frame_client_2_0212 = frame (4k, fill: [])
frame_client_2_0213 = frame (4k, fill: [])
frame_client_2_0214 = frame (4k, fill: [])
frame_client_2_0215 = frame (4k, fill: [])
frame_client_2_0216 = frame (4k, fill: [])
frame_client_2_0217 = frame (4k, fill: [])
frame_client_2_0218 = frame (4k, fill: [])
frame_client_2_0219 = frame (4k, fill: [])
frame_client_2_0220 = frame (4k, fill: [])
frame_client_2_0221 = frame (4k, fill: [])
frame_client_2_0222 = frame (4k, fill: [])
frame_client_2_0223 = frame (4k, fill: [])
frame_client_2_0224 = frame (4k, fill: [])
frame_client_2_0225 = frame (4k, fill: [])
frame_client_2_0226 = frame (4k, fill: [])
frame_client_2_0227 = frame (4k, fill: [])
frame_client_2_0228 = frame (4k, fill: [])
frame_client_2_0229 = frame (4k, fill: [])
frame_client_2_0230 = frame (4k, fill: [])
frame_client_2_0231 = frame (4k, fill: [])
frame_client_2_0232 = frame (4k, fill: [])
frame_client_2_0233 = frame (4k, fill: [])
frame_client_2_0234 = frame (4k, fill: [])
frame_client_2_0235 = frame (4k, fill: [])
frame_client_2_0236 = frame (4k, fill: [])
frame_client_2_0237 = frame (4k, fill: [])
frame_client_2_0238 = frame (4k, fill: [])
frame_client_2_0239 = frame (4k, fill: [])
frame_client_2_0240 = frame (4k, fill: [])
frame_client_2_0241 = frame (4k, fill: [])
frame_client_2_0242 = frame (4k, fill: [])
frame_client_2_0243 = frame (4k, fill: [])
frame_client_2_0244 = frame (4k, fill: [])
frame_client_2_0245 = frame (4k, fill: [])
frame_client_2_0246 = frame (4k, fill: [])
frame_client_2_0247 = frame (4k, fill: [])
frame_client_2_0248 = frame (4k, fill: [])
frame_client_2_0249 = frame (4k, fill: [])
frame_client_2_0250 = frame (4k, fill: [])
frame_client_2_0251 = frame (4k, fill: [])
frame_client_2_0252 = frame (4k, fill: [])
frame_client_2_0253 = frame (4k, fill: [])
frame_client_2_0254 = frame (4k, fill: [])
frame_client_2_0255 = frame (4k, fill: [])
frame_client_2_0256 = frame (4k, fill: [])
frame_client_2_0257 = frame (4k, fill: [])
frame_client_2_0258 = frame (4k, fill: [])
frame_client_2_0259 = frame (4k, fill: [])
frame_client_2_0260 = frame (4k, fill: [])
frame_client_2_0261 = frame (4k, fill: [])
frame_client_2_0262 = frame (4k, fill: [])
frame_client_2_0263 = frame (4k, fill: [])
frame_client_2_0264 = frame (4k, fill: [])
frame_client_2_0265 = frame (4k, fill: [])
frame_client_2_0266 = frame (4k, fill: [])
frame_client_2_0267 = frame (4k, fill: [])
frame_client_2_0268 = frame (4k, fill: [])
frame_client_2_0269 = frame (4k, fill: [])
frame_client_2_0270 = frame (4k, fill: [])
frame_client_2_0271 = frame (4k, fill: [])
frame_client_2_0272 = frame (4k, fill: [])
frame_client_2_0273 = frame (4k, fill: [])
frame_client_2_0274 = frame (4k, fill: [])
frame_client_2_0275 = frame (4k, fill: [])
frame_client_2_0276 = frame (4k, fill: [])
frame_client_2_0277 = frame (4k, fill: [])
frame_client_2_0278 = frame (4k, fill: [])
frame_client_2_0279 = frame (4k, fill: [])
frame_client_2_0280 = frame (4k, fill: [])
frame_client_2_0281 = frame (4k, fill: [])
frame_client_2_0282 = frame (4k, fill: [])
frame_client_2_0283 = frame (4k, fill: [])
frame_client_2_0284 = frame (4k, fill: [])
frame_client_2_0285 = frame (4k, fill: [])
frame_client_2_0286 = frame (4k, fill: [])
frame_client_2_0287 = frame (4k, fill: [])
frame_client_2_0288 = frame (4k, fill: [])
frame_client_2_0289 = frame (4k, fill: [])
frame_client_2_0290 = frame (4k, fill: [])
frame_client_2_0291 = frame (4k, fill: [])
frame_client_2_0292 = frame (4k, fill: [])
frame_client_2_0293 = frame (4k, fill: [])
frame_client_2_0294 = frame (4k, fill: [])
frame_client_2_0295 = frame (4k, fill: [])
frame_client_2_0296 = frame (4k, fill: [])
frame_client_2_0297 = frame (4k, fill: [])
frame_client_2_0298 = frame (4k, fill: [])
frame_client_2_0299 = frame (4k, fill: [])
frame_client_2_0300 = frame (4k, fill: [])
frame_client_2_0301 = frame (4k, fill: [])
frame_client_2_0302 = frame (4k, fill: [])
frame_client_2_0303 = frame (4k, fill: [])
frame_client_2_0304 = frame (4k, fill: [])
frame_client_2_0305 = frame (4k, fill: [])
frame_server_0000 = frame (4k, fill: [{0 548 CDL_FrameFill_FileData "server" 0}])
frame_server_0001 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "server" 4096}])
frame_server_0002 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "server" 8192}])
frame_server_0003 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "server" 12288}])
frame_server_0004 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "server" 16384}])
frame_server_0005 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "server" 20480}])
frame_server_0006 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "server" 24576}])
frame_server_0007 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "server" 28672}])
frame_server_0008 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "server" 32768}])
frame_server_0009 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "server" 36864}])
frame_server_0010 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "server" 40960}])
frame_server_0011 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "server" 45056}])
frame_server_0012 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "server" 49152}])
frame_server_0013 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "server" 53248}])
frame_server_0014 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "server" 57344}])
frame_server_0015 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "server" 61440}])
frame_server_0016 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "server" 65536}])
frame_server_0017 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "server" 69632}])
frame_server_0018 = frame (4k, fill: [{0 544 CDL_FrameFill_FileData "server" 73728}])
frame_server_0019 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "server" 77824}])
frame_server_0020 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "server" 81920}])
frame_server_0021 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "server" 86016}])
frame_server_0022 = frame (4k, fill: [{0 3056 CDL_FrameFill_FileData "server" 90112}])
frame_server_0023 = frame (4k, fill: [{4040 56 CDL_FrameFill_FileData "server" 94152}])
frame_server_0024 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "server" 94208}])
frame_server_0025 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "server" 98304}])
frame_server_0043 = frame (4k, fill: [{0 8 CDL_FrameFill_FileData "server" 172032}])
frame_server_0044 = frame (4k, fill: [])
frame_server_0045 = frame (4k, fill: [])
frame_server_0046 = frame (4k, fill: [])
frame_server_0047 = frame (4k, fill: [])
frame_server_0048 = frame (4k, fill: [])
frame_server_0049 = frame (4k, fill: [])
frame_server_0050 = frame (4k, fill: [])
frame_server_0051 = frame (4k, fill: [])
frame_server_0052 = frame (4k, fill: [])
frame_server_0053 = frame (4k, fill: [])
frame_server_0054 = frame (4k, fill: [])
frame_server_0055 = frame (4k, fill: [])
frame_server_0056 = frame (4k, fill: [])
frame_server_0057 = frame (4k, fill: [])
frame_server_0058 = frame (4k, fill: [])
frame_server_0059 = frame (4k, fill: [])
frame_server_0060 = frame (4k, fill: [])
frame_server_0061 = frame (4k, fill: [])
frame_server_0062 = frame (4k, fill: [])
frame_server_0063 = frame (4k, fill: [])
frame_server_0064 = frame (4k, fill: [])
frame_server_0065 = frame (4k, fill: [])
frame_server_0066 = frame (4k, fill: [])
frame_server_0067 = frame (4k, fill: [])
frame_server_0068 = frame (4k, fill: [])
frame_server_0069 = frame (4k, fill: [])
frame_server_0070 = frame (4k, fill: [])
frame_server_0071 = frame (4k, fill: [])
frame_server_0072 = frame (4k, fill: [])
frame_server_0073 = frame (4k, fill: [])
frame_server_0074 = frame (4k, fill: [])
frame_server_0075 = frame (4k, fill: [])
frame_server_0076 = frame (4k, fill: [])
frame_server_0077 = frame (4k, fill: [])
frame_server_0078 = frame (4k, fill: [])
frame_server_0079 = frame (4k, fill: [])
frame_server_0080 = frame (4k, fill: [])
frame_server_0081 = frame (4k, fill: [])
frame_server_0082 = frame (4k, fill: [])
frame_server_0083 = frame (4k, fill: [])
frame_server_0084 = frame (4k, fill: [])
frame_server_0085 = frame (4k, fill: [])
frame_server_0086 = frame (4k, fill: [])
frame_server_0087 = frame (4k, fill: [])
frame_server_0088 = frame (4k, fill: [])
frame_server_0089 = frame (4k, fill: [])
frame_server_0090 = frame (4k, fill: [])
frame_server_0091 = frame (4k, fill: [])
frame_server_0092 = frame (4k, fill: [])
frame_server_0093 = frame (4k, fill: [])
frame_server_0094 = frame (4k, fill: [])
frame_server_0095 = frame (4k, fill: [])
frame_server_0096 = frame (4k, fill: [])
frame_server_0097 = frame (4k, fill: [])
frame_server_0098 = frame (4k, fill: [])
frame_server_0099 = frame (4k, fill: [])
frame_server_0100 = frame (4k, fill: [])
frame_server_0101 = frame (4k, fill: [])
frame_server_0102 = frame (4k, fill: [])
frame_server_0103 = frame (4k, fill: [])
frame_server_0104 = frame (4k, fill: [])
frame_server_0105 = frame (4k, fill: [])
frame_server_0106 = frame (4k, fill: [])
frame_server_0107 = frame (4k, fill: [])
frame_server_0108 = frame (4k, fill: [])
frame_server_0109 = frame (4k, fill: [])
frame_server_0110 = frame (4k, fill: [])
frame_server_0111 = frame (4k, fill: [])
frame_server_0112 = frame (4k, fill: [])
frame_server_0113 = frame (4k, fill: [])
frame_server_0114 = frame (4k, fill: [])
frame_server_0115 = frame (4k, fill: [])
frame_server_0116 = frame (4k, fill: [])
frame_server_0117 = frame (4k, fill: [])
frame_server_0118 = frame (4k, fill: [])
frame_server_0119 = frame (4k, fill: [])
frame_server_0120 = frame (4k, fill: [])
frame_server_0121 = frame (4k, fill: [])
frame_server_0122 = frame (4k, fill: [])
frame_server_0123 = frame (4k, fill: [])
frame_server_0124 = frame (4k, fill: [])
frame_server_0125 = frame (4k, fill: [])
frame_server_0126 = frame (4k, fill: [])
frame_server_0127 = frame (4k, fill: [])
frame_server_0128 = frame (4k, fill: [])
frame_server_0129 = frame (4k, fill: [])
frame_server_0130 = frame (4k, fill: [])
frame_server_0131 = frame (4k, fill: [])
frame_server_0132 = frame (4k, fill: [])
frame_server_0133 = frame (4k, fill: [])
frame_server_0134 = frame (4k, fill: [])
frame_server_0135 = frame (4k, fill: [])
frame_server_0136 = frame (4k, fill: [])
frame_server_0137 = frame (4k, fill: [])
frame_server_0138 = frame (4k, fill: [])
frame_server_0139 = frame (4k, fill: [])
frame_server_0140 = frame (4k, fill: [])
frame_server_0141 = frame (4k, fill: [])
frame_server_0142 = frame (4k, fill: [])
frame_server_0143 = frame (4k, fill: [])
frame_server_0144 = frame (4k, fill: [])
frame_server_0145 = frame (4k, fill: [])
frame_server_0146 = frame (4k, fill: [])
frame_server_0147 = frame (4k, fill: [])
frame_server_0148 = frame (4k, fill: [])
frame_server_0149 = frame (4k, fill: [])
frame_server_0150 = frame (4k, fill: [])
frame_server_0151 = frame (4k, fill: [])
frame_server_0152 = frame (4k, fill: [])
frame_server_0153 = frame (4k, fill: [])
frame_server_0154 = frame (4k, fill: [])
frame_server_0155 = frame (4k, fill: [])
frame_server_0156 = frame (4k, fill: [])
frame_server_0157 = frame (4k, fill: [])
frame_server_0158 = frame (4k, fill: [])
frame_server_0159 = frame (4k, fill: [])
frame_server_0160 = frame (4k, fill: [])
frame_server_0161 = frame (4k, fill: [])
frame_server_0162 = frame (4k, fill: [])
frame_server_0163 = frame (4k, fill: [])
frame_server_0164 = frame (4k, fill: [])
frame_server_0165 = frame (4k, fill: [])
frame_server_0166 = frame (4k, fill: [])
frame_server_0167 = frame (4k, fill: [])
frame_server_0168 = frame (4k, fill: [])
frame_server_0169 = frame (4k, fill: [])
frame_server_0170 = frame (4k, fill: [])
frame_server_0171 = frame (4k, fill: [])
frame_server_0172 = frame (4k, fill: [])
frame_server_0173 = frame (4k, fill: [])
frame_server_0174 = frame (4k, fill: [])
frame_server_0175 = frame (4k, fill: [])
frame_server_0176 = frame (4k, fill: [])
frame_server_0177 = frame (4k, fill: [])
frame_server_0178 = frame (4k, fill: [])
frame_server_0179 = frame (4k, fill: [])
frame_server_0180 = frame (4k, fill: [])
frame_server_0181 = frame (4k, fill: [])
frame_server_0182 = frame (4k, fill: [])
frame_server_0183 = frame (4k, fill: [])
frame_server_0184 = frame (4k, fill: [])
frame_server_0185 = frame (4k, fill: [])
frame_server_0186 = frame (4k, fill: [])
frame_server_0187 = frame (4k, fill: [])
frame_server_0188 = frame (4k, fill: [])
frame_server_0189 = frame (4k, fill: [])
frame_server_0190 = frame (4k, fill: [])
frame_server_0191 = frame (4k, fill: [])
frame_server_0192 = frame (4k, fill: [])
frame_server_0193 = frame (4k, fill: [])
frame_server_0194 = frame (4k, fill: [])
frame_server_0195 = frame (4k, fill: [])
frame_server_0196 = frame (4k, fill: [])
frame_server_0197 = frame (4k, fill: [])
frame_server_0198 = frame (4k, fill: [])
frame_server_0199 = frame (4k, fill: [])
frame_server_0200 = frame (4k, fill: [])
frame_server_0201 = frame (4k, fill: [])
frame_server_0202 = frame (4k, fill: [])
frame_server_0203 = frame (4k, fill: [])
frame_server_0204 = frame (4k, fill: [])
frame_server_0205 = frame (4k, fill: [])
frame_server_0206 = frame (4k, fill: [])
frame_server_0207 = frame (4k, fill: [])
frame_server_0208 = frame (4k, fill: [])
frame_server_0209 = frame (4k, fill: [])
frame_server_0210 = frame (4k, fill: [])
frame_server_0211 = frame (4k, fill: [])
frame_server_0212 = frame (4k, fill: [])
frame_server_0213 = frame (4k, fill: [])
frame_server_0214 = frame (4k, fill: [])
frame_server_0215 = frame (4k, fill: [])
frame_server_0216 = frame (4k, fill: [])
frame_server_0217 = frame (4k, fill: [])
frame_server_0218 = frame (4k, fill: [])
frame_server_0219 = frame (4k, fill: [])
frame_server_0220 = frame (4k, fill: [])
frame_server_0221 = frame (4k, fill: [])
frame_server_0222 = frame (4k, fill: [])
frame_server_0223 = frame (4k, fill: [])
frame_server_0224 = frame (4k, fill: [])
frame_server_0225 = frame (4k, fill: [])
frame_server_0226 = frame (4k, fill: [])
frame_server_0227 = frame (4k, fill: [])
frame_server_0228 = frame (4k, fill: [])
frame_server_0229 = frame (4k, fill: [])
frame_server_0230 = frame (4k, fill: [])
frame_server_0231 = frame (4k, fill: [])
frame_server_0232 = frame (4k, fill: [])
frame_server_0233 = frame (4k, fill: [])
frame_server_0234 = frame (4k, fill: [])
frame_server_0235 = frame (4k, fill: [])
frame_server_0236 = frame (4k, fill: [])
frame_server_0237 = frame (4k, fill: [])
frame_server_0238 = frame (4k, fill: [])
frame_server_0239 = frame (4k, fill: [])
frame_server_0240 = frame (4k, fill: [])
frame_server_0241 = frame (4k, fill: [])
frame_server_0242 = frame (4k, fill: [])
frame_server_0243 = frame (4k, fill: [])
frame_server_0244 = frame (4k, fill: [])
frame_server_0245 = frame (4k, fill: [])
frame_server_0246 = frame (4k, fill: [])
frame_server_0247 = frame (4k, fill: [])
frame_server_0248 = frame (4k, fill: [])
frame_server_0249 = frame (4k, fill: [])
frame_server_0250 = frame (4k, fill: [])
frame_server_0251 = frame (4k, fill: [])
frame_server_0252 = frame (4k, fill: [])
frame_server_0253 = frame (4k, fill: [])
frame_server_0254 = frame (4k, fill: [])
frame_server_0255 = frame (4k, fill: [])
frame_server_0256 = frame (4k, fill: [])
frame_server_0257 = frame (4k, fill: [])
frame_server_0258 = frame (4k, fill: [])
frame_server_0259 = frame (4k, fill: [])
frame_server_0260 = frame (4k, fill: [])
frame_server_0261 = frame (4k, fill: [])
frame_server_0262 = frame (4k, fill: [])
frame_server_0263 = frame (4k, fill: [])
frame_server_0264 = frame (4k, fill: [])
frame_server_0265 = frame (4k, fill: [])
frame_server_0266 = frame (4k, fill: [])
frame_server_0267 = frame (4k, fill: [])
frame_server_0268 = frame (4k, fill: [])
frame_server_0269 = frame (4k, fill: [])
frame_server_0270 = frame (4k, fill: [])
frame_server_0271 = frame (4k, fill: [])
frame_server_0272 = frame (4k, fill: [])
frame_server_0273 = frame (4k, fill: [])
frame_server_0274 = frame (4k, fill: [])
frame_server_0275 = frame (4k, fill: [])
frame_server_0276 = frame (4k, fill: [])
frame_server_0277 = frame (4k, fill: [])
frame_server_0278 = frame (4k, fill: [])
frame_server_0279 = frame (4k, fill: [])
frame_server_0280 = frame (4k, fill: [])
frame_server_0281 = frame (4k, fill: [])
frame_server_0282 = frame (4k, fill: [])
frame_server_0283 = frame (4k, fill: [])
frame_server_0284 = frame (4k, fill: [])
frame_server_0285 = frame (4k, fill: [])
frame_server_0286 = frame (4k, fill: [])
frame_server_0287 = frame (4k, fill: [])
frame_server_0288 = frame (4k, fill: [])
frame_server_0289 = frame (4k, fill: [])
frame_server_0290 = frame (4k, fill: [])
frame_server_0291 = frame (4k, fill: [])
frame_server_0292 = frame (4k, fill: [])
frame_server_0293 = frame (4k, fill: [])
frame_server_0294 = frame (4k, fill: [])
frame_server_0295 = frame (4k, fill: [])
frame_server_0296 = frame (4k, fill: [])
frame_server_0297 = frame (4k, fill: [])
frame_server_0298 = frame (4k, fill: [])
frame_server_0299 = frame (4k, fill: [])
frame_server_0300 = frame (4k, fill: [])
frame_server_0301 = frame (4k, fill: [])
frame_server_0302 = frame (4k, fill: [])
frame_server_0303 = frame (4k, fill: [])
frame_server_0304 = frame (4k, fill: [])
frame_server_0305 = frame (4k, fill: [])
frame_server_0306 = frame (4k, fill: [])
ipc_client_1_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_1" 163840}])
ipc_client_2_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_2" 163840}])
ipc_server_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "server" 167936}])
pd_client_1_0001 = pd
pd_client_2_0001 = pd
pd_server_0001 = pd
pdpt_client_1_0000 = pdpt
pdpt_client_2_0000 = pdpt
pdpt_server_0000 = pdpt
pt_client_1_0002 = pt
pt_client_2_0002 = pt
pt_server_0002 = pt
stack_0_client_1_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_1" 98304}])
stack_0_client_2_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_2" 98304}])
stack_0_server_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "server" 102400}])
stack_10_client_1_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_1" 139264}])
stack_10_client_2_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_2" 139264}])
stack_10_server_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "server" 143360}])
stack_11_client_1_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_1" 143360}])
stack_11_client_2_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_2" 143360}])
stack_11_server_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "server" 147456}])
stack_12_client_1_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_1" 147456}])
stack_12_client_2_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_2" 147456}])
stack_12_server_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "server" 151552}])
stack_13_client_1_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_1" 151552}])
stack_13_client_2_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_2" 151552}])
stack_13_server_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "server" 155648}])
stack_14_client_1_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_1" 155648}])
stack_14_client_2_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_2" 155648}])
stack_14_server_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "server" 159744}])
stack_15_client_1_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_1" 159744}])
stack_15_client_2_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_2" 159744}])
stack_15_server_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "server" 163840}])
stack_1_client_1_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_1" 102400}])
stack_1_client_2_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_2" 102400}])
stack_1_server_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "server" 106496}])
stack_2_client_1_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_1" 106496}])
stack_2_client_2_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_2" 106496}])
stack_2_server_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "server" 110592}])
stack_3_client_1_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_1" 110592}])
stack_3_client_2_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_2" 110592}])
stack_3_server_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "server" 114688}])
stack_4_client_1_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_1" 114688}])
stack_4_client_2_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_2" 114688}])
stack_4_server_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "server" 118784}])
stack_5_client_1_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_1" 118784}])
stack_5_client_2_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_2" 118784}])
stack_5_server_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "server" 122880}])
stack_6_client_1_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_1" 122880}])
stack_6_client_2_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_2" 122880}])
stack_6_server_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "server" 126976}])
stack_7_client_1_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_1" 126976}])
stack_7_client_2_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_2" 126976}])
stack_7_server_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "server" 131072}])
stack_8_client_1_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_1" 131072}])
stack_8_client_2_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_2" 131072}])
stack_8_server_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "server" 135168}])
stack_9_client_1_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_1" 135168}])
stack_9_client_2_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "client_2" 135168}])
stack_9_server_obj = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "server" 139264}])
tcb_client_1 = tcb (addr: 0x429000,ip: 0x40103a,sp: 0x41a000,prio: 254,max_prio: 254,affinity: 0,init: [0, 0, 0, 0, 2, 4288600, 1, 0, 0, 32, 4209171, 0, 0])
tcb_client_2 = tcb (addr: 0x429000,ip: 0x40103a,sp: 0x41a000,prio: 254,max_prio: 254,affinity: 0,init: [0, 0, 0, 0, 2, 4288608, 1, 0, 0, 32, 4209171, 0, 0])
tcb_server = tcb (addr: 0x42a000,ip: 0x40103a,sp: 0x41b000,prio: 254,max_prio: 254,affinity: 0,init: [0, 0, 0, 0, 2, 4292640, 1, 0, 0, 32, 4211426, 0, 0])
vspace_client_1 = pml4
vspace_client_2 = pml4
vspace_server = pml4
}

caps {
cnode_client_1 {
0x1: endpoint (RWG)
0x2: cnode_client_1 (guard: 0, guard_size: 61)
0x4: tcb_client_1
}
cnode_client_2 {
0x1: endpoint (RWG)
0x2: cnode_client_2 (guard: 0, guard_size: 61)
0x4: tcb_client_2
}
cnode_server {
0x1: endpoint (RWG)
0x2: cnode_server (guard: 0, guard_size: 61)
0x4: tcb_server
}
pd_client_1_0001 {
0x2: pt_client_1_0002
}
pd_client_2_0001 {
0x2: pt_client_2_0002
}
pd_server_0001 {
0x2: pt_server_0002
}
pdpt_client_1_0000 {
0x0: pd_client_1_0001
}
pdpt_client_2_0000 {
0x0: pd_client_2_0001
}
pdpt_server_0000 {
0x0: pd_server_0001
}
pt_client_1_0002 {
0x0: frame_client_1_0000 (R)
0x1: frame_client_1_0001 (RX)
0x2: frame_client_1_0002 (RX)
0x3: frame_client_1_0003 (RX)
0x4: frame_client_1_0004 (RX)
0x5: frame_client_1_0005 (RX)
0x6: frame_client_1_0006 (RX)
0x7: frame_client_1_0007 (RX)
0x8: frame_client_1_0008 (RX)
0x9: frame_client_1_0009 (RX)
0xa: frame_client_1_0010 (RX)
0xb: frame_client_1_0011 (RX)
0xc: frame_client_1_0012 (RX)
0xd: frame_client_1_0013 (RX)
0xe: frame_client_1_0014 (RX)
0xf: frame_client_1_0015 (RX)
0x10: frame_client_1_0016 (RX)
0x11: frame_client_1_0017 (RX)
0x12: frame_client_1_0018 (R)
0x13: frame_client_1_0019 (R)
0x14: frame_client_1_0020 (R)
0x15: frame_client_1_0021 (R)
0x16: frame_client_1_0022 (RW)
0x17: frame_client_1_0023 (RW)
0x18: frame_client_1_0024 (RW)
0x19: stack_0_client_1_obj (RW)
0x1a: stack_1_client_1_obj (RW)
0x1b: stack_2_client_1_obj (RW)
0x1c: stack_3_client_1_obj (RW)
0x1d: stack_4_client_1_obj (RW)
0x1e: stack_5_client_1_obj (RW)
0x1f: stack_6_client_1_obj (RW)
0x20: stack_7_client_1_obj (RW)
0x21: stack_8_client_1_obj (RW)
0x22: stack_9_client_1_obj (RW)
0x23: stack_10_client_1_obj (RW)
0x24: stack_11_client_1_obj (RW)
0x25: stack_12_client_1_obj (RW)
0x26: stack_13_client_1_obj (RW)
0x27: stack_14_client_1_obj (RW)
0x28: stack_15_client_1_obj (RW)
0x29: ipc_client_1_obj (RW)
0x2a: frame_client_1_0042 (RW)
0x2b: frame_client_1_0043 (RW)
0x2c: frame_client_1_0044 (RW)
0x2d: frame_client_1_0045 (RW)
0x2e: frame_client_1_0046 (RW)
0x2f: frame_client_1_0047 (RW)
0x30: frame_client_1_0048 (RW)
0x31: frame_client_1_0049 (RW)
0x32: frame_client_1_0050 (RW)
0x33: frame_client_1_0051 (RW)
0x34: frame_client_1_0052 (RW)
0x35: frame_client_1_0053 (RW)
0x36: frame_client_1_0054 (RW)
0x37: frame_client_1_0055 (RW)
0x38: frame_client_1_0056 (RW)
0x39: frame_client_1_0057 (RW)
0x3a: frame_client_1_0058 (RW)
0x3b: frame_client_1_0059 (RW)
0x3c: frame_client_1_0060 (RW)
0x3d: frame_client_1_0061 (RW)
0x3e: frame_client_1_0062 (RW)
0x3f: frame_client_1_0063 (RW)
0x40: frame_client_1_0064 (RW)
0x41: frame_client_1_0065 (RW)
0x42: frame_client_1_0066 (RW)
0x43: frame_client_1_0067 (RW)
0x44: frame_client_1_0068 (RW)
0x45: frame_client_1_0069 (RW)
0x46: frame_client_1_0070 (RW)
0x47: frame_client_1_0071 (RW)
0x48: frame_client_1_0072 (RW)
0x49: frame_client_1_0073 (RW)
0x4a: frame_client_1_0074 (RW)
0x4b: frame_client_1_0075 (RW)
0x4c: frame_client_1_0076 (RW)
0x4d: frame_client_1_0077 (RW)
0x4e: frame_client_1_0078 (RW)
0x4f: frame_client_1_0079 (RW)
0x50: frame_client_1_0080 (RW)
0x51: frame_client_1_0081 (RW)
0x52: frame_client_1_0082 (RW)
0x53: frame_client_1_0083 (RW)
0x54: frame_client_1_0084 (RW)
0x55: frame_client_1_0085 (RW)
0x56: frame_client_1_0086 (RW)
0x57: frame_client_1_0087 (RW)
0x58: frame_client_1_0088 (RW)
0x59: frame_client_1_0089 (RW)
0x5a: frame_client_1_0090 (RW)
0x5b: frame_client_1_0091 (RW)
0x5c: frame_client_1_0092 (RW)
0x5d: frame_client_1_0093 (RW)
0x5e: frame_client_1_0094 (RW)
0x5f: frame_client_1_0095 (RW)
0x60: frame_client_1_0096 (RW)
0x61: frame_client_1_0097 (RW)
0x62: frame_client_1_0098 (RW)
0x63: frame_client_1_0099 (RW)
0x64: frame_client_1_0100 (RW)
0x65: frame_client_1_0101 (RW)
0x66: frame_client_1_0102 (RW)
0x67: frame_client_1_0103 (RW)
0x68: frame_client_1_0104 (RW)
0x69: frame_client_1_0105 (RW)
0x6a: frame_client_1_0106 (RW)
0x6b: frame_client_1_0107 (RW)
0x6c: frame_client_1_0108 (RW)
0x6d: frame_client_1_0109 (RW)
0x6e: frame_client_1_0110 (RW)
0x6f: frame_client_1_0111 (RW)
0x70: frame_client_1_0112 (RW)
0x71: frame_client_1_0113 (RW)
0x72: frame_client_1_0114 (RW)
0x73: frame_client_1_0115 (RW)
0x74: frame_client_1_0116 (RW)
0x75: frame_client_1_0117 (RW)
0x76: frame_client_1_0118 (RW)
0x77: frame_client_1_0119 (RW)
0x78: frame_client_1_0120 (RW)
0x79: frame_client_1_0121 (RW)
0x7a: frame_client_1_0122 (RW)
0x7b: frame_client_1_0123 (RW)
0x7c: frame_client_1_0124 (RW)
0x7d: frame_client_1_0125 (RW)
0x7e: frame_client_1_0126 (RW)
0x7f: frame_client_1_0127 (RW)
0x80: frame_client_1_0128 (RW)
0x81: frame_client_1_0129 (RW)
0x82: frame_client_1_0130 (RW)
0x83: frame_client_1_0131 (RW)
0x84: frame_client_1_0132 (RW)
0x85: frame_client_1_0133 (RW)
0x86: frame_client_1_0134 (RW)
0x87: frame_client_1_0135 (RW)
0x88: frame_client_1_0136 (RW)
0x89: frame_client_1_0137 (RW)
0x8a: frame_client_1_0138 (RW)
0x8b: frame_client_1_0139 (RW)
0x8c: frame_client_1_0140 (RW)
0x8d: frame_client_1_0141 (RW)
0x8e: frame_client_1_0142 (RW)
0x8f: frame_client_1_0143 (RW)
0x90: frame_client_1_0144 (RW)
0x91: frame_client_1_0145 (RW)
0x92: frame_client_1_0146 (RW)
0x93: frame_client_1_0147 (RW)
0x94: frame_client_1_0148 (RW)
0x95: frame_client_1_0149 (RW)
0x96: frame_client_1_0150 (RW)
0x97: frame_client_1_0151 (RW)
0x98: frame_client_1_0152 (RW)
0x99: frame_client_1_0153 (RW)
0x9a: frame_client_1_0154 (RW)
0x9b: frame_client_1_0155 (RW)
0x9c: frame_client_1_0156 (RW)
0x9d: frame_client_1_0157 (RW)
0x9e: frame_client_1_0158 (RW)
0x9f: frame_client_1_0159 (RW)
0xa0: frame_client_1_0160 (RW)
0xa1: frame_client_1_0161 (RW)
0xa2: frame_client_1_0162 (RW)
0xa3: frame_client_1_0163 (RW)
0xa4: frame_client_1_0164 (RW)
0xa5: frame_client_1_0165 (RW)
0xa6: frame_client_1_0166 (RW)
0xa7: frame_client_1_0167 (RW)
0xa8: frame_client_1_0168 (RW)
0xa9: frame_client_1_0169 (RW)
0xaa: frame_client_1_0170 (RW)
0xab: frame_client_1_0171 (RW)
0xac: frame_client_1_0172 (RW)
0xad: frame_client_1_0173 (RW)
0xae: frame_client_1_0174 (RW)
0xaf: frame_client_1_0175 (RW)
0xb0: frame_client_1_0176 (RW)
0xb1: frame_client_1_0177 (RW)
0xb2: frame_client_1_0178 (RW)
0xb3: frame_client_1_0179 (RW)
0xb4: frame_client_1_0180 (RW)
0xb5: frame_client_1_0181 (RW)
0xb6: frame_client_1_0182 (RW)
0xb7: frame_client_1_0183 (RW)
0xb8: frame_client_1_0184 (RW)
0xb9: frame_client_1_0185 (RW)
0xba: frame_client_1_0186 (RW)
0xbb: frame_client_1_0187 (RW)
0xbc: frame_client_1_0188 (RW)
0xbd: frame_client_1_0189 (RW)
0xbe: frame_client_1_0190 (RW)
0xbf: frame_client_1_0191 (RW)
0xc0: frame_client_1_0192 (RW)
0xc1: frame_client_1_0193 (RW)
0xc2: frame_client_1_0194 (RW)
0xc3: frame_client_1_0195 (RW)
0xc4: frame_client_1_0196 (RW)
0xc5: frame_client_1_0197 (RW)
0xc6: frame_client_1_0198 (RW)
0xc7: frame_client_1_0199 (RW)
0xc8: frame_client_1_0200 (RW)
0xc9: frame_client_1_0201 (RW)
0xca: frame_client_1_0202 (RW)
0xcb: frame_client_1_0203 (RW)
0xcc: frame_client_1_0204 (RW)
0xcd: frame_client_1_0205 (RW)
0xce: frame_client_1_0206 (RW)
0xcf: frame_client_1_0207 (RW)
0xd0: frame_client_1_0208 (RW)
0xd1: frame_client_1_0209 (RW)
0xd2: frame_client_1_0210 (RW)
0xd3: frame_client_1_0211 (RW)
0xd4: frame_client_1_0212 (RW)
0xd5: frame_client_1_0213 (RW)
0xd6: frame_client_1_0214 (RW)
0xd7: frame_client_1_0215 (RW)
0xd8: frame_client_1_0216 (RW)
0xd9: frame_client_1_0217 (RW)
0xda: frame_client_1_0218 (RW)
0xdb: frame_client_1_0219 (RW)
0xdc: frame_client_1_0220 (RW)
0xdd: frame_client_1_0221 (RW)
0xde: frame_client_1_0222 (RW)
0xdf: frame_client_1_0223 (RW)
0xe0: frame_client_1_0224 (RW)
0xe1: frame_client_1_0225 (RW)
0xe2: frame_client_1_0226 (RW)
0xe3: frame_client_1_0227 (RW)
0xe4: frame_client_1_0228 (RW)
0xe5: frame_client_1_0229 (RW)
0xe6: frame_client_1_0230 (RW)
0xe7: frame_client_1_0231 (RW)
0xe8: frame_client_1_0232 (RW)
0xe9: frame_client_1_0233 (RW)
0xea: frame_client_1_0234 (RW)
0xeb: frame_client_1_0235 (RW)
0xec: frame_client_1_0236 (RW)
0xed: frame_client_1_0237 (RW)
0xee: frame_client_1_0238 (RW)
0xef: frame_client_1_0239 (RW)
0xf0: frame_client_1_0240 (RW)
0xf1: frame_client_1_0241 (RW)
0xf2: frame_client_1_0242 (RW)
0xf3: frame_client_1_0243 (RW)
0xf4: frame_client_1_0244 (RW)
0xf5: frame_client_1_0245 (RW)
0xf6: frame_client_1_0246 (RW)
0xf7: frame_client_1_0247 (RW)
0xf8: frame_client_1_0248 (RW)
0xf9: frame_client_1_0249 (RW)
0xfa: frame_client_1_0250 (RW)
0xfb: frame_client_1_0251 (RW)
0xfc: frame_client_1_0252 (RW)
0xfd: frame_client_1_0253 (RW)
0xfe: frame_client_1_0254 (RW)
0xff: frame_client_1_0255 (RW)
0x100: frame_client_1_0256 (RW)
0x101: frame_client_1_0257 (RW)
0x102: frame_client_1_0258 (RW)
0x103: frame_client_1_0259 (RW)
0x104: frame_client_1_0260 (RW)
0x105: frame_client_1_0261 (RW)
0x106: frame_client_1_0262 (RW)
0x107: frame_client_1_0263 (RW)
0x108: frame_client_1_0264 (RW)
0x109: frame_client_1_0265 (RW)
0x10a: frame_client_1_0266 (RW)
0x10b: frame_client_1_0267 (RW)
0x10c: frame_client_1_0268 (RW)
0x10d: frame_client_1_0269 (RW)
0x10e: frame_client_1_0270 (RW)
0x10f: frame_client_1_0271 (RW)
0x110: frame_client_1_0272 (RW)
0x111: frame_client_1_0273 (RW)
0x112: frame_client_1_0274 (RW)
0x113: frame_client_1_0275 (RW)
0x114: frame_client_1_0276 (RW)
0x115: frame_client_1_0277 (RW)
0x116: frame_client_1_0278 (RW)
0x117: frame_client_1_0279 (RW)
0x118: frame_client_1_0280 (RW)
0x119: frame_client_1_0281 (RW)
0x11a: frame_client_1_0282 (RW)
0x11b: frame_client_1_0283 (RW)
0x11c: frame_client_1_0284 (RW)
0x11d: frame_client_1_0285 (RW)
0x11e: frame_client_1_0286 (RW)
0x11f: frame_client_1_0287 (RW)
0x120: frame_client_1_0288 (RW)
0x121: frame_client_1_0289 (RW)
0x122: frame_client_1_0290 (RW)
0x123: frame_client_1_0291 (RW)
0x124: frame_client_1_0292 (RW)
0x125: frame_client_1_0293 (RW)
0x126: frame_client_1_0294 (RW)
0x127: frame_client_1_0295 (RW)
0x128: frame_client_1_0296 (RW)
0x129: frame_client_1_0297 (RW)
0x12a: frame_client_1_0298 (RW)
0x12b: frame_client_1_0299 (RW)
0x12c: frame_client_1_0300 (RW)
0x12d: frame_client_1_0301 (RW)
0x12e: frame_client_1_0302 (RW)
0x12f: frame_client_1_0303 (RW)
0x130: frame_client_1_0304 (RW)
0x131: frame_client_1_0305 (RW)
}
pt_client_2_0002 {
0x0: frame_client_2_0000 (R)
0x1: frame_client_2_0001 (RX)
0x2: frame_client_2_0002 (RX)
0x3: frame_client_2_0003 (RX)
0x4: frame_client_2_0004 (RX)
0x5: frame_client_2_0005 (RX)
0x6: frame_client_2_0006 (RX)
0x7: frame_client_2_0007 (RX)
0x8: frame_client_2_0008 (RX)
0x9: frame_client_2_0009 (RX)
0xa: frame_client_2_0010 (RX)
0xb: frame_client_2_0011 (RX)
0xc: frame_client_2_0012 (RX)
0xd: frame_client_2_0013 (RX)
0xe: frame_client_2_0014 (RX)
0xf: frame_client_2_0015 (RX)
0x10: frame_client_2_0016 (RX)
0x11: frame_client_2_0017 (RX)
0x12: frame_client_2_0018 (R)
0x13: frame_client_2_0019 (R)
0x14: frame_client_2_0020 (R)
0x15: frame_client_2_0021 (R)
0x16: frame_client_2_0022 (RW)
0x17: frame_client_2_0023 (RW)
0x18: frame_client_2_0024 (RW)
0x19: stack_0_client_2_obj (RW)
0x1a: stack_1_client_2_obj (RW)
0x1b: stack_2_client_2_obj (RW)
0x1c: stack_3_client_2_obj (RW)
0x1d: stack_4_client_2_obj (RW)
0x1e: stack_5_client_2_obj (RW)
0x1f: stack_6_client_2_obj (RW)
0x20: stack_7_client_2_obj (RW)
0x21: stack_8_client_2_obj (RW)
0x22: stack_9_client_2_obj (RW)
0x23: stack_10_client_2_obj (RW)
0x24: stack_11_client_2_obj (RW)
0x25: stack_12_client_2_obj (RW)
0x26: stack_13_client_2_obj (RW)
0x27: stack_14_client_2_obj (RW)
0x28: stack_15_client_2_obj (RW)
0x29: ipc_client_2_obj (RW)
0x2a: frame_client_2_0042 (RW)
0x2b: frame_client_2_0043 (RW)
0x2c: frame_client_2_0044 (RW)
0x2d: frame_client_2_0045 (RW)
0x2e: frame_client_2_0046 (RW)
0x2f: frame_client_2_0047 (RW)
0x30: frame_client_2_0048 (RW)
0x31: frame_client_2_0049 (RW)
0x32: frame_client_2_0050 (RW)
0x33: frame_client_2_0051 (RW)
0x34: frame_client_2_0052 (RW)
0x35: frame_client_2_0053 (RW)
0x36: frame_client_2_0054 (RW)
0x37: frame_client_2_0055 (RW)
0x38: frame_client_2_0056 (RW)
0x39: frame_client_2_0057 (RW)
0x3a: frame_client_2_0058 (RW)
0x3b: frame_client_2_0059 (RW)
0x3c: frame_client_2_0060 (RW)
0x3d: frame_client_2_0061 (RW)
0x3e: frame_client_2_0062 (RW)
0x3f: frame_client_2_0063 (RW)
0x40: frame_client_2_0064 (RW)
0x41: frame_client_2_0065 (RW)
0x42: frame_client_2_0066 (RW)
0x43: frame_client_2_0067 (RW)
0x44: frame_client_2_0068 (RW)
0x45: frame_client_2_0069 (RW)
0x46: frame_client_2_0070 (RW)
0x47: frame_client_2_0071 (RW)
0x48: frame_client_2_0072 (RW)
0x49: frame_client_2_0073 (RW)
0x4a: frame_client_2_0074 (RW)
0x4b: frame_client_2_0075 (RW)
0x4c: frame_client_2_0076 (RW)
0x4d: frame_client_2_0077 (RW)
0x4e: frame_client_2_0078 (RW)
0x4f: frame_client_2_0079 (RW)
0x50: frame_client_2_0080 (RW)
0x51: frame_client_2_0081 (RW)
0x52: frame_client_2_0082 (RW)
0x53: frame_client_2_0083 (RW)
0x54: frame_client_2_0084 (RW)
0x55: frame_client_2_0085 (RW)
0x56: frame_client_2_0086 (RW)
0x57: frame_client_2_0087 (RW)
0x58: frame_client_2_0088 (RW)
0x59: frame_client_2_0089 (RW)
0x5a: frame_client_2_0090 (RW)
0x5b: frame_client_2_0091 (RW)
0x5c: frame_client_2_0092 (RW)
0x5d: frame_client_2_0093 (RW)
0x5e: frame_client_2_0094 (RW)
0x5f: frame_client_2_0095 (RW)
0x60: frame_client_2_0096 (RW)
0x61: frame_client_2_0097 (RW)
0x62: frame_client_2_0098 (RW)
0x63: frame_client_2_0099 (RW)
0x64: frame_client_2_0100 (RW)
0x65: frame_client_2_0101 (RW)
0x66: frame_client_2_0102 (RW)
0x67: frame_client_2_0103 (RW)
0x68: frame_client_2_0104 (RW)
0x69: frame_client_2_0105 (RW)
0x6a: frame_client_2_0106 (RW)
0x6b: frame_client_2_0107 (RW)
0x6c: frame_client_2_0108 (RW)
0x6d: frame_client_2_0109 (RW)
0x6e: frame_client_2_0110 (RW)
0x6f: frame_client_2_0111 (RW)
0x70: frame_client_2_0112 (RW)
0x71: frame_client_2_0113 (RW)
0x72: frame_client_2_0114 (RW)
0x73: frame_client_2_0115 (RW)
0x74: frame_client_2_0116 (RW)
0x75: frame_client_2_0117 (RW)
0x76: frame_client_2_0118 (RW)
0x77: frame_client_2_0119 (RW)
0x78: frame_client_2_0120 (RW)
0x79: frame_client_2_0121 (RW)
0x7a: frame_client_2_0122 (RW)
0x7b: frame_client_2_0123 (RW)
0x7c: frame_client_2_0124 (RW)
0x7d: frame_client_2_0125 (RW)
0x7e: frame_client_2_0126 (RW)
0x7f: frame_client_2_0127 (RW)
0x80: frame_client_2_0128 (RW)
0x81: frame_client_2_0129 (RW)
0x82: frame_client_2_0130 (RW)
0x83: frame_client_2_0131 (RW)
0x84: frame_client_2_0132 (RW)
0x85: frame_client_2_0133 (RW)
0x86: frame_client_2_0134 (RW)
0x87: frame_client_2_0135 (RW)
0x88: frame_client_2_0136 (RW)
0x89: frame_client_2_0137 (RW)
0x8a: frame_client_2_0138 (RW)
0x8b: frame_client_2_0139 (RW)
0x8c: frame_client_2_0140 (RW)
0x8d: frame_client_2_0141 (RW)
0x8e: frame_client_2_0142 (RW)
0x8f: frame_client_2_0143 (RW)
0x90: frame_client_2_0144 (RW)
0x91: frame_client_2_0145 (RW)
0x92: frame_client_2_0146 (RW)
0x93: frame_client_2_0147 (RW)
0x94: frame_client_2_0148 (RW)
0x95: frame_client_2_0149 (RW)
0x96: frame_client_2_0150 (RW)
0x97: frame_client_2_0151 (RW)
0x98: frame_client_2_0152 (RW)
0x99: frame_client_2_0153 (RW)
0x9a: frame_client_2_0154 (RW)
0x9b: frame_client_2_0155 (RW)
0x9c: frame_client_2_0156 (RW)
0x9d: frame_client_2_0157 (RW)
0x9e: frame_client_2_0158 (RW)
0x9f: frame_client_2_0159 (RW)
0xa0: frame_client_2_0160 (RW)
0xa1: frame_client_2_0161 (RW)
0xa2: frame_client_2_0162 (RW)
0xa3: frame_client_2_0163 (RW)
0xa4: frame_client_2_0164 (RW)
0xa5: frame_client_2_0165 (RW)
0xa6: frame_client_2_0166 (RW)
0xa7: frame_client_2_0167 (RW)
0xa8: frame_client_2_0168 (RW)
0xa9: frame_client_2_0169 (RW)
0xaa: frame_client_2_0170 (RW)
0xab: frame_client_2_0171 (RW)
0xac: frame_client_2_0172 (RW)
0xad: frame_client_2_0173 (RW)
0xae: frame_client_2_0174 (RW)
0xaf: frame_client_2_0175 (RW)
0xb0: frame_client_2_0176 (RW)
0xb1: frame_client_2_0177 (RW)
0xb2: frame_client_2_0178 (RW)
0xb3: frame_client_2_0179 (RW)
0xb4: frame_client_2_0180 (RW)
0xb5: frame_client_2_0181 (RW)
0xb6: frame_client_2_0182 (RW)
0xb7: frame_client_2_0183 (RW)
0xb8: frame_client_2_0184 (RW)
0xb9: frame_client_2_0185 (RW)
0xba: frame_client_2_0186 (RW)
0xbb: frame_client_2_0187 (RW)
0xbc: frame_client_2_0188 (RW)
0xbd: frame_client_2_0189 (RW)
0xbe: frame_client_2_0190 (RW)
0xbf: frame_client_2_0191 (RW)
0xc0: frame_client_2_0192 (RW)
0xc1: frame_client_2_0193 (RW)
0xc2: frame_client_2_0194 (RW)
0xc3: frame_client_2_0195 (RW)
0xc4: frame_client_2_0196 (RW)
0xc5: frame_client_2_0197 (RW)
0xc6: frame_client_2_0198 (RW)
0xc7: frame_client_2_0199 (RW)
0xc8: frame_client_2_0200 (RW)
0xc9: frame_client_2_0201 (RW)
0xca: frame_client_2_0202 (RW)
0xcb: frame_client_2_0203 (RW)
0xcc: frame_client_2_0204 (RW)
0xcd: frame_client_2_0205 (RW)
0xce: frame_client_2_0206 (RW)
0xcf: frame_client_2_0207 (RW)
0xd0: frame_client_2_0208 (RW)
0xd1: frame_client_2_0209 (RW)
0xd2: frame_client_2_0210 (RW)
0xd3: frame_client_2_0211 (RW)
0xd4: frame_client_2_0212 (RW)
0xd5: frame_client_2_0213 (RW)
0xd6: frame_client_2_0214 (RW)
0xd7: frame_client_2_0215 (RW)
0xd8: frame_client_2_0216 (RW)
0xd9: frame_client_2_0217 (RW)
0xda: frame_client_2_0218 (RW)
0xdb: frame_client_2_0219 (RW)
0xdc: frame_client_2_0220 (RW)
0xdd: frame_client_2_0221 (RW)
0xde: frame_client_2_0222 (RW)
0xdf: frame_client_2_0223 (RW)
0xe0: frame_client_2_0224 (RW)
0xe1: frame_client_2_0225 (RW)
0xe2: frame_client_2_0226 (RW)
0xe3: frame_client_2_0227 (RW)
0xe4: frame_client_2_0228 (RW)
0xe5: frame_client_2_0229 (RW)
0xe6: frame_client_2_0230 (RW)
0xe7: frame_client_2_0231 (RW)
0xe8: frame_client_2_0232 (RW)
0xe9: frame_client_2_0233 (RW)
0xea: frame_client_2_0234 (RW)
0xeb: frame_client_2_0235 (RW)
0xec: frame_client_2_0236 (RW)
0xed: frame_client_2_0237 (RW)
0xee: frame_client_2_0238 (RW)
0xef: frame_client_2_0239 (RW)
0xf0: frame_client_2_0240 (RW)
0xf1: frame_client_2_0241 (RW)
0xf2: frame_client_2_0242 (RW)
0xf3: frame_client_2_0243 (RW)
0xf4: frame_client_2_0244 (RW)
0xf5: frame_client_2_0245 (RW)
0xf6: frame_client_2_0246 (RW)
0xf7: frame_client_2_0247 (RW)
0xf8: frame_client_2_0248 (RW)
0xf9: frame_client_2_0249 (RW)
0xfa: frame_client_2_0250 (RW)
0xfb: frame_client_2_0251 (RW)
0xfc: frame_client_2_0252 (RW)
0xfd: frame_client_2_0253 (RW)
0xfe: frame_client_2_0254 (RW)
0xff: frame_client_2_0255 (RW)
0x100: frame_client_2_0256 (RW)
0x101: frame_client_2_0257 (RW)
0x102: frame_client_2_0258 (RW)
0x103: frame_client_2_0259 (RW)
0x104: frame_client_2_0260 (RW)
0x105: frame_client_2_0261 (RW)
0x106: frame_client_2_0262 (RW)
0x107: frame_client_2_0263 (RW)
0x108: frame_client_2_0264 (RW)
0x109: frame_client_2_0265 (RW)
0x10a: frame_client_2_0266 (RW)
0x10b: frame_client_2_0267 (RW)
0x10c: frame_client_2_0268 (RW)
0x10d: frame_client_2_0269 (RW)
0x10e: frame_client_2_0270 (RW)
0x10f: frame_client_2_0271 (RW)
0x110: frame_client_2_0272 (RW)
0x111: frame_client_2_0273 (RW)
0x112: frame_client_2_0274 (RW)
0x113: frame_client_2_0275 (RW)
0x114: frame_client_2_0276 (RW)
0x115: frame_client_2_0277 (RW)
0x116: frame_client_2_0278 (RW)
0x117: frame_client_2_0279 (RW)
0x118: frame_client_2_0280 (RW)
0x119: frame_client_2_0281 (RW)
0x11a: frame_client_2_0282 (RW)
0x11b: frame_client_2_0283 (RW)
0x11c: frame_client_2_0284 (RW)
0x11d: frame_client_2_0285 (RW)
0x11e: frame_client_2_0286 (RW)
0x11f: frame_client_2_0287 (RW)
0x120: frame_client_2_0288 (RW)
0x121: frame_client_2_0289 (RW)
0x122: frame_client_2_0290 (RW)
0x123: frame_client_2_0291 (RW)
0x124: frame_client_2_0292 (RW)
0x125: frame_client_2_0293 (RW)
0x126: frame_client_2_0294 (RW)
0x127: frame_client_2_0295 (RW)
0x128: frame_client_2_0296 (RW)
0x129: frame_client_2_0297 (RW)
0x12a: frame_client_2_0298 (RW)
0x12b: frame_client_2_0299 (RW)
0x12c: frame_client_2_0300 (RW)
0x12d: frame_client_2_0301 (RW)
0x12e: frame_client_2_0302 (RW)
0x12f: frame_client_2_0303 (RW)
0x130: frame_client_2_0304 (RW)
0x131: frame_client_2_0305 (RW)
}
pt_server_0002 {
0x0: frame_server_0000 (R)
0x1: frame_server_0001 (RX)
0x2: frame_server_0002 (RX)
0x3: frame_server_0003 (RX)
0x4: frame_server_0004 (RX)
0x5: frame_server_0005 (RX)
0x6: frame_server_0006 (RX)
0x7: frame_server_0007 (RX)
0x8: frame_server_0008 (RX)
0x9: frame_server_0009 (RX)
0xa: frame_server_0010 (RX)
0xb: frame_server_0011 (RX)
0xc: frame_server_0012 (RX)
0xd: frame_server_0013 (RX)
0xe: frame_server_0014 (RX)
0xf: frame_server_0015 (RX)
0x10: frame_server_0016 (RX)
0x11: frame_server_0017 (RX)
0x12: frame_server_0018 (RX)
0x13: frame_server_0019 (R)
0x14: frame_server_0020 (R)
0x15: frame_server_0021 (R)
0x16: frame_server_0022 (R)
0x17: frame_server_0023 (RW)
0x18: frame_server_0024 (RW)
0x19: frame_server_0025 (RW)
0x1a: stack_0_server_obj (RW)
0x1b: stack_1_server_obj (RW)
0x1c: stack_2_server_obj (RW)
0x1d: stack_3_server_obj (RW)
0x1e: stack_4_server_obj (RW)
0x1f: stack_5_server_obj (RW)
0x20: stack_6_server_obj (RW)
0x21: stack_7_server_obj (RW)
0x22: stack_8_server_obj (RW)
0x23: stack_9_server_obj (RW)
0x24: stack_10_server_obj (RW)
0x25: stack_11_server_obj (RW)
0x26: stack_12_server_obj (RW)
0x27: stack_13_server_obj (RW)
0x28: stack_14_server_obj (RW)
0x29: stack_15_server_obj (RW)
0x2a: ipc_server_obj (RW)
0x2b: frame_server_0043 (RW)
0x2c: frame_server_0044 (RW)
0x2d: frame_server_0045 (RW)
0x2e: frame_server_0046 (RW)
0x2f: frame_server_0047 (RW)
0x30: frame_server_0048 (RW)
0x31: frame_server_0049 (RW)
0x32: frame_server_0050 (RW)
0x33: frame_server_0051 (RW)
0x34: frame_server_0052 (RW)
0x35: frame_server_0053 (RW)
0x36: frame_server_0054 (RW)
0x37: frame_server_0055 (RW)
0x38: frame_server_0056 (RW)
0x39: frame_server_0057 (RW)
0x3a: frame_server_0058 (RW)
0x3b: frame_server_0059 (RW)
0x3c: frame_server_0060 (RW)
0x3d: frame_server_0061 (RW)
0x3e: frame_server_0062 (RW)
0x3f: frame_server_0063 (RW)
0x40: frame_server_0064 (RW)
0x41: frame_server_0065 (RW)
0x42: frame_server_0066 (RW)
0x43: frame_server_0067 (RW)
0x44: frame_server_0068 (RW)
0x45: frame_server_0069 (RW)
0x46: frame_server_0070 (RW)
0x47: frame_server_0071 (RW)
0x48: frame_server_0072 (RW)
0x49: frame_server_0073 (RW)
0x4a: frame_server_0074 (RW)
0x4b: frame_server_0075 (RW)
0x4c: frame_server_0076 (RW)
0x4d: frame_server_0077 (RW)
0x4e: frame_server_0078 (RW)
0x4f: frame_server_0079 (RW)
0x50: frame_server_0080 (RW)
0x51: frame_server_0081 (RW)
0x52: frame_server_0082 (RW)
0x53: frame_server_0083 (RW)
0x54: frame_server_0084 (RW)
0x55: frame_server_0085 (RW)
0x56: frame_server_0086 (RW)
0x57: frame_server_0087 (RW)
0x58: frame_server_0088 (RW)
0x59: frame_server_0089 (RW)
0x5a: frame_server_0090 (RW)
0x5b: frame_server_0091 (RW)
0x5c: frame_server_0092 (RW)
0x5d: frame_server_0093 (RW)
0x5e: frame_server_0094 (RW)
0x5f: frame_server_0095 (RW)
0x60: frame_server_0096 (RW)
0x61: frame_server_0097 (RW)
0x62: frame_server_0098 (RW)
0x63: frame_server_0099 (RW)
0x64: frame_server_0100 (RW)
0x65: frame_server_0101 (RW)
0x66: frame_server_0102 (RW)
0x67: frame_server_0103 (RW)
0x68: frame_server_0104 (RW)
0x69: frame_server_0105 (RW)
0x6a: frame_server_0106 (RW)
0x6b: frame_server_0107 (RW)
0x6c: frame_server_0108 (RW)
0x6d: frame_server_0109 (RW)
0x6e: frame_server_0110 (RW)
0x6f: frame_server_0111 (RW)
0x70: frame_server_0112 (RW)
0x71: frame_server_0113 (RW)
0x72: frame_server_0114 (RW)
0x73: frame_server_0115 (RW)
0x74: frame_server_0116 (RW)
0x75: frame_server_0117 (RW)
0x76: frame_server_0118 (RW)
0x77: frame_server_0119 (RW)
0x78: frame_server_0120 (RW)
0x79: frame_server_0121 (RW)
0x7a: frame_server_0122 (RW)
0x7b: frame_server_0123 (RW)
0x7c: frame_server_0124 (RW)
0x7d: frame_server_0125 (RW)
0x7e: frame_server_0126 (RW)
0x7f: frame_server_0127 (RW)
0x80: frame_server_0128 (RW)
0x81: frame_server_0129 (RW)
0x82: frame_server_0130 (RW)
0x83: frame_server_0131 (RW)
0x84: frame_server_0132 (RW)
0x85: frame_server_0133 (RW)
0x86: frame_server_0134 (RW)
0x87: frame_server_0135 (RW)
0x88: frame_server_0136 (RW)
0x89: frame_server_0137 (RW)
0x8a: frame_server_0138 (RW)
0x8b: frame_server_0139 (RW)
0x8c: frame_server_0140 (RW)
0x8d: frame_server_0141 (RW)
0x8e: frame_server_0142 (RW)
0x8f: frame_server_0143 (RW)
0x90: frame_server_0144 (RW)
0x91: frame_server_0145 (RW)
0x92: frame_server_0146 (RW)
0x93: frame_server_0147 (RW)
0x94: frame_server_0148 (RW)
0x95: frame_server_0149 (RW)
0x96: frame_server_0150 (RW)
0x97: frame_server_0151 (RW)
0x98: frame_server_0152 (RW)
0x99: frame_server_0153 (RW)
0x9a: frame_server_0154 (RW)
0x9b: frame_server_0155 (RW)
0x9c: frame_server_0156 (RW)
0x9d: frame_server_0157 (RW)
0x9e: frame_server_0158 (RW)
0x9f: frame_server_0159 (RW)
0xa0: frame_server_0160 (RW)
0xa1: frame_server_0161 (RW)
0xa2: frame_server_0162 (RW)
0xa3: frame_server_0163 (RW)
0xa4: frame_server_0164 (RW)
0xa5: frame_server_0165 (RW)
0xa6: frame_server_0166 (RW)
0xa7: frame_server_0167 (RW)
0xa8: frame_server_0168 (RW)
0xa9: frame_server_0169 (RW)
0xaa: frame_server_0170 (RW)
0xab: frame_server_0171 (RW)
0xac: frame_server_0172 (RW)
0xad: frame_server_0173 (RW)
0xae: frame_server_0174 (RW)
0xaf: frame_server_0175 (RW)
0xb0: frame_server_0176 (RW)
0xb1: frame_server_0177 (RW)
0xb2: frame_server_0178 (RW)
0xb3: frame_server_0179 (RW)
0xb4: frame_server_0180 (RW)
0xb5: frame_server_0181 (RW)
0xb6: frame_server_0182 (RW)
0xb7: frame_server_0183 (RW)
0xb8: frame_server_0184 (RW)
0xb9: frame_server_0185 (RW)
0xba: frame_server_0186 (RW)
0xbb: frame_server_0187 (RW)
0xbc: frame_server_0188 (RW)
0xbd: frame_server_0189 (RW)
0xbe: frame_server_0190 (RW)
0xbf: frame_server_0191 (RW)
0xc0: frame_server_0192 (RW)
0xc1: frame_server_0193 (RW)
0xc2: frame_server_0194 (RW)
0xc3: frame_server_0195 (RW)
0xc4: frame_server_0196 (RW)
0xc5: frame_server_0197 (RW)
0xc6: frame_server_0198 (RW)
0xc7: frame_server_0199 (RW)
0xc8: frame_server_0200 (RW)
0xc9: frame_server_0201 (RW)
0xca: frame_server_0202 (RW)
0xcb: frame_server_0203 (RW)
0xcc: frame_server_0204 (RW)
0xcd: frame_server_0205 (RW)
0xce: frame_server_0206 (RW)
0xcf: frame_server_0207 (RW)
0xd0: frame_server_0208 (RW)
0xd1: frame_server_0209 (RW)
0xd2: frame_server_0210 (RW)
0xd3: frame_server_0211 (RW)
0xd4: frame_server_0212 (RW)
0xd5: frame_server_0213 (RW)
0xd6: frame_server_0214 (RW)
0xd7: frame_server_0215 (RW)
0xd8: frame_server_0216 (RW)
0xd9: frame_server_0217 (RW)
0xda: frame_server_0218 (RW)
0xdb: frame_server_0219 (RW)
0xdc: frame_server_0220 (RW)
0xdd: frame_server_0221 (RW)
0xde: frame_server_0222 (RW)
0xdf: frame_server_0223 (RW)
0xe0: frame_server_0224 (RW)
0xe1: frame_server_0225 (RW)
0xe2: frame_server_0226 (RW)
0xe3: frame_server_0227 (RW)
0xe4: frame_server_0228 (RW)
0xe5: frame_server_0229 (RW)
0xe6: frame_server_0230 (RW)
0xe7: frame_server_0231 (RW)
0xe8: frame_server_0232 (RW)
0xe9: frame_server_0233 (RW)
0xea: frame_server_0234 (RW)
0xeb: frame_server_0235 (RW)
0xec: frame_server_0236 (RW)
0xed: frame_server_0237 (RW)
0xee: frame_server_0238 (RW)
0xef: frame_server_0239 (RW)
0xf0: frame_server_0240 (RW)
0xf1: frame_server_0241 (RW)
0xf2: frame_server_0242 (RW)
0xf3: frame_server_0243 (RW)
0xf4: frame_server_0244 (RW)
0xf5: frame_server_0245 (RW)
0xf6: frame_server_0246 (RW)
0xf7: frame_server_0247 (RW)
0xf8: frame_server_0248 (RW)
0xf9: frame_server_0249 (RW)
0xfa: frame_server_0250 (RW)
0xfb: frame_server_0251 (RW)
0xfc: frame_server_0252 (RW)
0xfd: frame_server_0253 (RW)
0xfe: frame_server_0254 (RW)
0xff: frame_server_0255 (RW)
0x100: frame_server_0256 (RW)
0x101: frame_server_0257 (RW)
0x102: frame_server_0258 (RW)
0x103: frame_server_0259 (RW)
0x104: frame_server_0260 (RW)
0x105: frame_server_0261 (RW)
0x106: frame_server_0262 (RW)
0x107: frame_server_0263 (RW)
0x108: frame_server_0264 (RW)
0x109: frame_server_0265 (RW)
0x10a: frame_server_0266 (RW)
0x10b: frame_server_0267 (RW)
0x10c: frame_server_0268 (RW)
0x10d: frame_server_0269 (RW)
0x10e: frame_server_0270 (RW)
0x10f: frame_server_0271 (RW)
0x110: frame_server_0272 (RW)
0x111: frame_server_0273 (RW)
0x112: frame_server_0274 (RW)
0x113: frame_server_0275 (RW)
0x114: frame_server_0276 (RW)
0x115: frame_server_0277 (RW)
0x116: frame_server_0278 (RW)
0x117: frame_server_0279 (RW)
0x118: frame_server_0280 (RW)
0x119: frame_server_0281 (RW)
0x11a: frame_server_0282 (RW)
0x11b: frame_server_0283 (RW)
0x11c: frame_server_0284 (RW)
0x11d: frame_server_0285 (RW)
0x11e: frame_server_0286 (RW)
0x11f: frame_server_0287 (RW)
0x120: frame_server_0288 (RW)
0x121: frame_server_0289 (RW)
0x122: frame_server_0290 (RW)
0x123: frame_server_0291 (RW)
0x124: frame_server_0292 (RW)
0x125: frame_server_0293 (RW)
0x126: frame_server_0294 (RW)
0x127: frame_server_0295 (RW)
0x128: frame_server_0296 (RW)
0x129: frame_server_0297 (RW)
0x12a: frame_server_0298 (RW)
0x12b: frame_server_0299 (RW)
0x12c: frame_server_0300 (RW)
0x12d: frame_server_0301 (RW)
0x12e: frame_server_0302 (RW)
0x12f: frame_server_0303 (RW)
0x130: frame_server_0304 (RW)
0x131: frame_server_0305 (RW)
0x132: frame_server_0306 (RW)
}
tcb_client_1 {
cspace: cnode_client_1 (guard: 0, guard_size: 61)
ipc_buffer_slot: ipc_client_1_obj (RW)
vspace: vspace_client_1
}
tcb_client_2 {
cspace: cnode_client_2 (guard: 0, guard_size: 61)
ipc_buffer_slot: ipc_client_2_obj (RW)
vspace: vspace_client_2
}
tcb_server {
cspace: cnode_server (guard: 0, guard_size: 61)
ipc_buffer_slot: ipc_server_obj (RW)
vspace: vspace_server
}
vspace_client_1 {
0x0: pdpt_client_1_0000
}
vspace_client_2 {
0x0: pdpt_client_2_0000
}
vspace_server {
0x0: pdpt_server_0000
}
}

irq maps {

}